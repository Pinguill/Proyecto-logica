-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Fri Jun 11 15:10:40 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY verificador IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        cont : IN STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
        outN : OUT STD_LOGIC;
        outP : OUT STD_LOGIC;
        outK : OUT STD_LOGIC;
        outTemp : OUT STD_LOGIC;
        outHum : OUT STD_LOGIC
    );
END verificador;

ARCHITECTURE BEHAVIOR OF verificador IS
    TYPE type_fstate IS (data,valN,valP,valK,valTemp,valHum);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,cont)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= data;
            outN <= '0';
            outP <= '0';
            outK <= '0';
            outTemp <= '0';
            outHum <= '0';
        ELSE
            outN <= '0';
            outP <= '0';
            outK <= '0';
            outTemp <= '0';
            outHum <= '0';
            CASE fstate IS
                WHEN data =>
                    IF ((cont(2 DOWNTO 0) = "000")) THEN
                        reg_fstate <= valN;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= data;
                    END IF;
                WHEN valN =>
                    IF ((cont(2 DOWNTO 0) = "001")) THEN
                        reg_fstate <= valP;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= valN;
                    END IF;

                    outN <= '1';
                WHEN valP =>
                    IF ((cont(2 DOWNTO 0) = "010")) THEN
                        reg_fstate <= valK;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= valP;
                    END IF;

                    outP <= '1';
                WHEN valK =>
                    IF ((cont(2 DOWNTO 0) = "011")) THEN
                        reg_fstate <= valTemp;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= valK;
                    END IF;

                    outK <= '1';
                WHEN valTemp =>
                    IF ((cont(2 DOWNTO 0) = "100")) THEN
                        reg_fstate <= valHum;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= valTemp;
                    END IF;

                    outTemp <= '1';
                WHEN valHum =>
                    reg_fstate <= data;

                    outHum <= '1';
                WHEN OTHERS => 
                    outN <= 'X';
                    outP <= 'X';
                    outK <= 'X';
                    outTemp <= 'X';
                    outHum <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
